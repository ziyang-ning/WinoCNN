
module data_controller ();

endmodule


module data_buffer ();

endmodule


module data_trans ();

endmodule


module data_top ();

endmodule

